`timescale 1ns / 1ps



module T_matris_rom(
    input wire clk_i,rst_i,rd_i, // senkron calismasi icin 
    input wire [5:0] addr_i, // romdaki adres bilgisi
    output reg [31:0] data_o
    );
    reg [31:0] ROM[0:63];  // 32 bitlik 2^6(64) satirlik bir rom
    
    initial begin
        ROM[0] = 32'b00111101111111111100101110010010; // 0.1249
        ROM[1] = 32'b00111110001101001111000011011000; // 0.1767
        ROM[2] = 32'b00111110001101001111000011011000;
        ROM[3] = 32'b00111110001101001111000011011000;
        ROM[4] = 32'b00111110001101001111000011011000;
        ROM[5] = 32'b00111110001101001111000011011000;
        ROM[6] = 32'b00111110001101001111000011011000;
        ROM[7] = 32'b00111110001101001111000011011000;
        ROM[8] = 32'b00111110001101001111000011011000; // 0,1767
        ROM[9] = 32'b00111110100000000000000000000000; // 0.25
        ROM[10] = 32'b00111110100000000000000000000000; 
        ROM[11] = 32'b00111110100000000000000000000000; 
        ROM[12] = 32'b00111110100000000000000000000000; 
        ROM[13] = 32'b00111110100000000000000000000000; 
        ROM[14] = 32'b00111110100000000000000000000000; 
        ROM[15] = 32'b00111110100000000000000000000000; 
        ROM[16] = 32'b00111110001101001111000011011000; // 0,1767
        ROM[17] = 32'b00111110100000000000000000000000; // 0.25
        ROM[18] = 32'b00111110100000000000000000000000; 
        ROM[19] = 32'b00111110100000000000000000000000; 
        ROM[20] = 32'b00111110100000000000000000000000; 
        ROM[21] = 32'b00111110100000000000000000000000; 
        ROM[22] = 32'b00111110100000000000000000000000; 
        ROM[23] = 32'b00111110100000000000000000000000; 
        ROM[24] = 32'b00111110001101001111000011011000; // 0,1767
        ROM[25] = 32'b00111110100000000000000000000000; // 0.25
        ROM[26] = 32'b00111110100000000000000000000000; 
        ROM[27] = 32'b00111110100000000000000000000000; 
        ROM[28] = 32'b00111110100000000000000000000000; 
        ROM[29] = 32'b00111110100000000000000000000000; 
        ROM[30] = 32'b00111110100000000000000000000000; 
        ROM[31] = 32'b00111110100000000000000000000000; 
        ROM[32] = 32'b00111110001101001111000011011000; // 0,1767
        ROM[33] = 32'b00111110100000000000000000000000; // 0.25
        ROM[34] = 32'b00111110100000000000000000000000; 
        ROM[35] = 32'b00111110100000000000000000000000; 
        ROM[36] = 32'b00111110100000000000000000000000; 
        ROM[37] = 32'b00111110100000000000000000000000; 
        ROM[38] = 32'b00111110100000000000000000000000; 
        ROM[39] = 32'b00111110100000000000000000000000; 
        ROM[40] = 32'b00111110001101001111000011011000; // 0,1767
        ROM[41] = 32'b00111110100000000000000000000000; // 0.25
        ROM[42] = 32'b00111110100000000000000000000000; 
        ROM[43] = 32'b00111110100000000000000000000000; 
        ROM[44] = 32'b00111110100000000000000000000000; 
        ROM[45] = 32'b00111110100000000000000000000000; 
        ROM[46] = 32'b00111110100000000000000000000000; 
        ROM[47] = 32'b00111110100000000000000000000000; 
        ROM[48] = 32'b00111110001101001111000011011000; // 0,1767
        ROM[49] = 32'b00111110100000000000000000000000; // 0.25
        ROM[50] = 32'b00111110100000000000000000000000; 
        ROM[51] = 32'b00111110100000000000000000000000; 
        ROM[52] = 32'b00111110100000000000000000000000; 
        ROM[53] = 32'b00111110100000000000000000000000; 
        ROM[54] = 32'b00111110100000000000000000000000; 
        ROM[55] = 32'b00111110100000000000000000000000; 
        ROM[56] = 32'b00111110001101001111000011011000; // 0,1767
        ROM[57] = 32'b00111110100000000000000000000000; // 0.25
        ROM[58] = 32'b00111110100000000000000000000000; 
        ROM[59] = 32'b00111110100000000000000000000000; 
        ROM[60] = 32'b00111110100000000000000000000000; 
        ROM[61] = 32'b00111110100000000000000000000000; 
        ROM[62] = 32'b00111110100000000000000000000000; 
        ROM[63] = 32'b00111110100000000000000000000000; 
     end
                
        always @(posedge clk_i) begin
            if(rst_i)begin
            end else begin
               if(rd_i == 1)begin
                   data_o <= ROM[addr_i];
               end else begin
               end
            end
        end
        

endmodule
