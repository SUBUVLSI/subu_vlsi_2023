`timescale 1ns / 1ps

module kuantalama_rom(
    input wire clk_i,rst_i,rd_i,  // senkron calismasi icin 
    input wire [5:0] addr_i, // romdaki adres bilgisi 
    output reg signed [10:0] data_o
    );
    reg signed [10:0] ROM[0:63];  // 11 bitlik, 2^6(64) satirlik bir işaretli rom
    
    initial begin
        ROM[0] = 11'b00000010000; // 16
        ROM[1] = 11'b00000001011; // 11
        ROM[2] = 11'b00000001010; // 10
        ROM[3] = 11'b00000010000; // 16
        ROM[4] = 11'b00000011000; // 24
        ROM[5] = 11'b00000101000; // 40
        ROM[6] = 11'b00000110011; // 51
        ROM[7] = 11'b00000111101; // 61
        ROM[8] = 11'b00000001100; // 12
        ROM[9] = 11'b00000001100; // 12
        ROM[10] = 11'b00000001110; // 14
        ROM[11] = 11'b00000010011; // 19
        ROM[12] = 11'b00000011010; // 26
        ROM[13] = 11'b00000111010; // 58
        ROM[14] = 11'b00000111100; // 60
        ROM[15] = 11'b00000110111; // 55
        ROM[16] = 11'b00000001110; // 14
        ROM[17] = 11'b00000001101; // 13
        ROM[18] = 11'b00000010000; // 16 
        ROM[19] = 11'b00000011000; // 24  
        ROM[20] = 11'b00000101000; // 40  
        ROM[21] = 11'b00000111001; // 57
        ROM[22] = 11'b00001000101; // 69
        ROM[23] = 11'b00000111000; // 56
        ROM[24] = 11'b00000001110; // 14
        ROM[25] = 11'b00000010001; // 17
        ROM[26] = 11'b00000010110; // 22
        ROM[27] = 11'b00000011101; // 29
        ROM[28] = 11'b00000110011; // 51
        ROM[29] = 11'b00001010111; // 87
        ROM[30] = 11'b00001010000; // 80
        ROM[31] = 11'b00000111110; // 62
        ROM[32] = 11'b00000010010; // 18
        ROM[33] = 11'b00000010110; // 22 
        ROM[34] = 11'b00000100101; // 37
        ROM[35] = 11'b00000111000; // 56 
        ROM[36] = 11'b00001000100; // 68
        ROM[37] = 11'b00001101101; // 109
        ROM[38] = 11'b00001100111; // 103
        ROM[39] = 11'b00001001101; // 77
        ROM[40] = 11'b00000011000; // 24 
        ROM[41] = 11'b00000100011; // 35
        ROM[42] = 11'b00000110111; // 55
        ROM[43] = 11'b00001000000; // 64
        ROM[44] = 11'b00001010001; // 81
        ROM[45] = 11'b00001101000; // 104
        ROM[46] = 11'b00001110001; // 113
        ROM[47] = 11'b00001011100; // 92
        ROM[48] = 11'b00000110001; // 49
        ROM[49] = 11'b00001000000; // 64
        ROM[50] = 11'b00001001110; // 78
        ROM[51] = 11'b00001010111; // 87
        ROM[52] = 11'b00001100111; // 103
        ROM[53] = 11'b00001111001; // 121
        ROM[54] = 11'b00001111000; // 120
        ROM[55] = 11'b00001100101; // 101
        ROM[56] = 11'b00001001000; // 72
        ROM[57] = 11'b00001011100; // 92
        ROM[58] = 11'b00001011111; // 95
        ROM[59] = 11'b00001100010; // 98
        ROM[60] = 11'b00001110000; // 112
        ROM[61] = 11'b00001100100; // 100
        ROM[62] = 11'b00001100111; // 103
        ROM[63] = 11'b00001100011; // 99
     end
                
     always @(posedge clk_i) begin
         if(rst_i)begin
         end else begin
            if(rd_i == 1)begin
                data_o <= ROM[addr_i];
            end else begin
            end
         end
     end
        
endmodule
