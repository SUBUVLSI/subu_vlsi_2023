`timescale 1ns / 1ps

module kuantalama_rom(
    input wire clk_i,  // senkron calismasi icin 
    input wire [12:0] addr_i, // romdaki adres bilgisi 
    output reg signed [32:0] data_o
    );
    reg [31:0] ROM[0:5];  // 32 bitlik, 2^6(64) satirlik bir rom
    
    initial begin
        ROM[0] = 32'b01000001100000000000000000000000; // 16
        ROM[1] = 32'b01000001001100000000000000000000; // 11
        ROM[2] = 32'b01000001001000000000000000000000; // 10
        ROM[3] = 32'b01000001100000000000000000000000; // 16
        ROM[4] = 32'b01000001110000000000000000000000; // 24
        ROM[5] = 32'b01000010001000000000000000000000; // 40
        ROM[6] = 32'b01000010010011000000000000000000; // 51
        ROM[7] = 32'b01000010011101000000000000000000; // 61
        ROM[8] = 32'b01000001010000000000000000000000; // 12
        ROM[9] = 32'b01000001010000000000000000000000; // 12
        ROM[10] = 32'b01000001011000000000000000000000; // 14
        ROM[11] = 32'b01000001100110000000000000000000; // 19
        ROM[12] = 32'b01000001110100000000000000000000; // 26
        ROM[13] = 32'b01000010011010000000000000000000; // 58
        ROM[14] = 32'b01000010011100000000000000000000; // 60
        ROM[15] = 32'b01000010010111000000000000000000; // 55
        ROM[16] = 32'b01000001011000000000000000000000; // 14
        ROM[17] = 32'b01000001010100000000000000000000; // 13
        ROM[18] = 32'b01000001100000000000000000000000; // 16 
        ROM[19] = 32'b01000001110000000000000000000000; // 24  
        ROM[20] = 32'b01000010001000000000000000000000; // 40  
        ROM[21] = 32'b01000010011001000000000000000000; // 57
        ROM[22] = 32'b01000010100010100000000000000000; // 69
        ROM[23] = 32'b01000010011000000000000000000000; // 56
        ROM[24] = 32'b01000001011000000000000000000000; // 14
        ROM[25] = 32'b01000001100010000000000000000000; // 17
        ROM[26] = 32'b01000001101100000000000000000000; // 22
        ROM[27] = 32'b01000001111010000000000000000000; // 29
        ROM[28] = 32'b01000010010011000000000000000000; // 51
        ROM[29] = 32'b01000010101011100000000000000000; // 87
        ROM[30] = 32'b01000010101000000000000000000000; // 80
        ROM[31] = 32'b01000010011110000000000000000000; // 62
        ROM[32] = 32'b01000001100100000000000000000000; // 18
        ROM[33] = 32'b01000001101100000000000000000000; // 22 
        ROM[34] = 32'b01000010000101000000000000000000; // 37
        ROM[35] = 32'b01000010011000000000000000000000; // 56 
        ROM[36] = 32'b01000010100010000000000000000000; // 68
        ROM[37] = 32'b01000010110110100000000000000000; // 109
        ROM[38] = 32'b01000010110011100000000000000000; // 103
        ROM[39] = 32'b01000010100110100000000000000000; // 77
        ROM[40] = 32'b01000001110000000000000000000000; // 24 
        ROM[41] = 32'b01000010000011000000000000000000; // 35
        ROM[42] = 32'b01000010010111000000000000000000; // 55
        ROM[43] = 32'b01000010100000000000000000000000; // 64
        ROM[44] = 32'b01000010101000100000000000000000; // 81
        ROM[45] = 32'b01000010110100000000000000000000; // 104
        ROM[46] = 32'b01000010111000100000000000000000; // 113
        ROM[47] = 32'b01000010101110000000000000000000; // 92
        ROM[48] = 32'b01000010010001000000000000000000; // 49
        ROM[49] = 32'b01000010100000000000000000000000; // 64
        ROM[50] = 32'b01000010100111000000000000000000; // 78
        ROM[51] = 32'b01000010101011100000000000000000; // 87
        ROM[52] = 32'b01000010110011100000000000000000; // 103
        ROM[53] = 32'b01000010111100100000000000000000; // 121
        ROM[54] = 32'b01000010111100000000000000000000; // 120
        ROM[55] = 32'b01000010110010100000000000000000; // 101
        ROM[56] = 32'b01000010100100000000000000000000; // 72
        ROM[57] = 32'b01000010101110000000000000000000; // 92
        ROM[58] = 32'b01000010101111100000000000000000; // 95
        ROM[59] = 32'b01000010110001000000000000000000; // 98
        ROM[60] = 32'b01000010111000000000000000000000; // 112
        ROM[61] = 32'b01000010110010000000000000000000; // 100
        ROM[62] = 32'b01000010110011100000000000000000; // 103
        ROM[63] = 32'b01000010110001100000000000000000; // 99
     end
                
        always @(posedge clk_i) begin
            data_o = ROM[addr_i];
        end
        

endmodule
